// projeto1.v

// Generated using ACDS version 13.1 162 at 2018.09.16.11:16:11

`timescale 1 ps / 1 ps
module projeto1 (
		input  wire  clk_clk,                                    //                                 clk.clk
		input  wire  reset_reset_n,                              //                               reset.reset_n
		input  wire  botaosubir_external_connection_export,      //      botaosubir_external_connection.export
		input  wire  botaodescer_external_connection_export,     //     botaodescer_external_connection.export
		input  wire  botaoselecionar_external_connection_export, // botaoselecionar_external_connection.export
		input  wire  botaovoltar_external_connection_export,     //     botaovoltar_external_connection.export
		output wire  ledopcao1_external_connection_export,       //       ledopcao1_external_connection.export
		output wire  ledopcao2_external_connection_export,       //       ledopcao2_external_connection.export
		output wire  ledopcao3_external_connection_export,       //       ledopcao3_external_connection.export
		output wire  ledopcao4_external_connection_export,       //       ledopcao4_external_connection.export
		output wire  ledopcao5_external_connection_export        //       ledopcao5_external_connection.export
	);

	wire   [1:0] mm_interconnect_0_botaodescer_s1_address;                     // mm_interconnect_0:botaoDescer_s1_address -> botaoDescer:address
	wire  [31:0] mm_interconnect_0_botaodescer_s1_readdata;                    // botaoDescer:readdata -> mm_interconnect_0:botaoDescer_s1_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [15:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire  [31:0] mm_interconnect_0_ledopcao4_s1_writedata;                     // mm_interconnect_0:ledOpcao4_s1_writedata -> ledOpcao4:writedata
	wire   [1:0] mm_interconnect_0_ledopcao4_s1_address;                       // mm_interconnect_0:ledOpcao4_s1_address -> ledOpcao4:address
	wire         mm_interconnect_0_ledopcao4_s1_chipselect;                    // mm_interconnect_0:ledOpcao4_s1_chipselect -> ledOpcao4:chipselect
	wire         mm_interconnect_0_ledopcao4_s1_write;                         // mm_interconnect_0:ledOpcao4_s1_write -> ledOpcao4:write_n
	wire  [31:0] mm_interconnect_0_ledopcao4_s1_readdata;                      // ledOpcao4:readdata -> mm_interconnect_0:ledOpcao4_s1_readdata
	wire   [1:0] mm_interconnect_0_botaoselecionar_s1_address;                 // mm_interconnect_0:botaoSelecionar_s1_address -> botaoSelecionar:address
	wire  [31:0] mm_interconnect_0_botaoselecionar_s1_readdata;                // botaoSelecionar:readdata -> mm_interconnect_0:botaoSelecionar_s1_readdata
	wire  [31:0] mm_interconnect_0_ledopcao1_s1_writedata;                     // mm_interconnect_0:ledOpcao1_s1_writedata -> ledOpcao1:writedata
	wire   [1:0] mm_interconnect_0_ledopcao1_s1_address;                       // mm_interconnect_0:ledOpcao1_s1_address -> ledOpcao1:address
	wire         mm_interconnect_0_ledopcao1_s1_chipselect;                    // mm_interconnect_0:ledOpcao1_s1_chipselect -> ledOpcao1:chipselect
	wire         mm_interconnect_0_ledopcao1_s1_write;                         // mm_interconnect_0:ledOpcao1_s1_write -> ledOpcao1:write_n
	wire  [31:0] mm_interconnect_0_ledopcao1_s1_readdata;                      // ledOpcao1:readdata -> mm_interconnect_0:ledOpcao1_s1_readdata
	wire  [31:0] mm_interconnect_0_ledopcao2_s1_writedata;                     // mm_interconnect_0:ledOpcao2_s1_writedata -> ledOpcao2:writedata
	wire   [1:0] mm_interconnect_0_ledopcao2_s1_address;                       // mm_interconnect_0:ledOpcao2_s1_address -> ledOpcao2:address
	wire         mm_interconnect_0_ledopcao2_s1_chipselect;                    // mm_interconnect_0:ledOpcao2_s1_chipselect -> ledOpcao2:chipselect
	wire         mm_interconnect_0_ledopcao2_s1_write;                         // mm_interconnect_0:ledOpcao2_s1_write -> ledOpcao2:write_n
	wire  [31:0] mm_interconnect_0_ledopcao2_s1_readdata;                      // ledOpcao2:readdata -> mm_interconnect_0:ledOpcao2_s1_readdata
	wire   [1:0] mm_interconnect_0_botaosubir_s1_address;                      // mm_interconnect_0:botaoSubir_s1_address -> botaoSubir:address
	wire  [31:0] mm_interconnect_0_botaosubir_s1_readdata;                     // botaoSubir:readdata -> mm_interconnect_0:botaoSubir_s1_readdata
	wire   [1:0] mm_interconnect_0_botaovoltar_s1_address;                     // mm_interconnect_0:botaoVoltar_s1_address -> botaoVoltar:address
	wire  [31:0] mm_interconnect_0_botaovoltar_s1_readdata;                    // botaoVoltar:readdata -> mm_interconnect_0:botaoVoltar_s1_readdata
	wire  [31:0] mm_interconnect_0_ledopcao5_s1_writedata;                     // mm_interconnect_0:ledOpcao5_s1_writedata -> ledOpcao5:writedata
	wire   [1:0] mm_interconnect_0_ledopcao5_s1_address;                       // mm_interconnect_0:ledOpcao5_s1_address -> ledOpcao5:address
	wire         mm_interconnect_0_ledopcao5_s1_chipselect;                    // mm_interconnect_0:ledOpcao5_s1_chipselect -> ledOpcao5:chipselect
	wire         mm_interconnect_0_ledopcao5_s1_write;                         // mm_interconnect_0:ledOpcao5_s1_write -> ledOpcao5:write_n
	wire  [31:0] mm_interconnect_0_ledopcao5_s1_readdata;                      // ledOpcao5:readdata -> mm_interconnect_0:ledOpcao5_s1_readdata
	wire  [31:0] mm_interconnect_0_ledopcao3_s1_writedata;                     // mm_interconnect_0:ledOpcao3_s1_writedata -> ledOpcao3:writedata
	wire   [1:0] mm_interconnect_0_ledopcao3_s1_address;                       // mm_interconnect_0:ledOpcao3_s1_address -> ledOpcao3:address
	wire         mm_interconnect_0_ledopcao3_s1_chipselect;                    // mm_interconnect_0:ledOpcao3_s1_chipselect -> ledOpcao3:chipselect
	wire         mm_interconnect_0_ledopcao3_s1_write;                         // mm_interconnect_0:ledOpcao3_s1_write -> ledOpcao3:write_n
	wire  [31:0] mm_interconnect_0_ledopcao3_s1_readdata;                      // ledOpcao3:readdata -> mm_interconnect_0:ledOpcao3_s1_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [15:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [botaoDescer:reset_n, botaoSelecionar:reset_n, botaoSubir:reset_n, botaoVoltar:reset_n, irq_mapper:reset, ledOpcao1:reset_n, ledOpcao2:reset_n, ledOpcao3:reset_n, ledOpcao4:reset_n, ledOpcao5:reset_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	projeto1_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                             //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	projeto1_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	projeto1_botaoSubir botaosubir (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_botaosubir_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botaosubir_s1_readdata), //                    .readdata
		.in_port  (botaosubir_external_connection_export)     // external_connection.export
	);

	projeto1_botaoSubir botaodescer (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_botaodescer_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botaodescer_s1_readdata), //                    .readdata
		.in_port  (botaodescer_external_connection_export)     // external_connection.export
	);

	projeto1_botaoSubir botaoselecionar (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_botaoselecionar_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botaoselecionar_s1_readdata), //                    .readdata
		.in_port  (botaoselecionar_external_connection_export)     // external_connection.export
	);

	projeto1_botaoSubir botaovoltar (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_botaovoltar_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botaovoltar_s1_readdata), //                    .readdata
		.in_port  (botaovoltar_external_connection_export)     // external_connection.export
	);

	projeto1_ledOpcao1 ledopcao1 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_ledopcao1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledopcao1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledopcao1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledopcao1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledopcao1_s1_readdata),   //                    .readdata
		.out_port   (ledopcao1_external_connection_export)       // external_connection.export
	);

	projeto1_ledOpcao1 ledopcao2 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_ledopcao2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledopcao2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledopcao2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledopcao2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledopcao2_s1_readdata),   //                    .readdata
		.out_port   (ledopcao2_external_connection_export)       // external_connection.export
	);

	projeto1_ledOpcao1 ledopcao3 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_ledopcao3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledopcao3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledopcao3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledopcao3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledopcao3_s1_readdata),   //                    .readdata
		.out_port   (ledopcao3_external_connection_export)       // external_connection.export
	);

	projeto1_ledOpcao1 ledopcao4 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_ledopcao4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledopcao4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledopcao4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledopcao4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledopcao4_s1_readdata),   //                    .readdata
		.out_port   (ledopcao4_external_connection_export)       // external_connection.export
	);

	projeto1_ledOpcao1 ledopcao5 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_ledopcao5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledopcao5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledopcao5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledopcao5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledopcao5_s1_readdata),   //                    .readdata
		.out_port   (ledopcao5_external_connection_export)       // external_connection.export
	);

	projeto1_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.botaoDescer_s1_address                           (mm_interconnect_0_botaodescer_s1_address),                     //                             botaoDescer_s1.address
		.botaoDescer_s1_readdata                          (mm_interconnect_0_botaodescer_s1_readdata),                    //                                           .readdata
		.botaoSelecionar_s1_address                       (mm_interconnect_0_botaoselecionar_s1_address),                 //                         botaoSelecionar_s1.address
		.botaoSelecionar_s1_readdata                      (mm_interconnect_0_botaoselecionar_s1_readdata),                //                                           .readdata
		.botaoSubir_s1_address                            (mm_interconnect_0_botaosubir_s1_address),                      //                              botaoSubir_s1.address
		.botaoSubir_s1_readdata                           (mm_interconnect_0_botaosubir_s1_readdata),                     //                                           .readdata
		.botaoVoltar_s1_address                           (mm_interconnect_0_botaovoltar_s1_address),                     //                             botaoVoltar_s1.address
		.botaoVoltar_s1_readdata                          (mm_interconnect_0_botaovoltar_s1_readdata),                    //                                           .readdata
		.ledOpcao1_s1_address                             (mm_interconnect_0_ledopcao1_s1_address),                       //                               ledOpcao1_s1.address
		.ledOpcao1_s1_write                               (mm_interconnect_0_ledopcao1_s1_write),                         //                                           .write
		.ledOpcao1_s1_readdata                            (mm_interconnect_0_ledopcao1_s1_readdata),                      //                                           .readdata
		.ledOpcao1_s1_writedata                           (mm_interconnect_0_ledopcao1_s1_writedata),                     //                                           .writedata
		.ledOpcao1_s1_chipselect                          (mm_interconnect_0_ledopcao1_s1_chipselect),                    //                                           .chipselect
		.ledOpcao2_s1_address                             (mm_interconnect_0_ledopcao2_s1_address),                       //                               ledOpcao2_s1.address
		.ledOpcao2_s1_write                               (mm_interconnect_0_ledopcao2_s1_write),                         //                                           .write
		.ledOpcao2_s1_readdata                            (mm_interconnect_0_ledopcao2_s1_readdata),                      //                                           .readdata
		.ledOpcao2_s1_writedata                           (mm_interconnect_0_ledopcao2_s1_writedata),                     //                                           .writedata
		.ledOpcao2_s1_chipselect                          (mm_interconnect_0_ledopcao2_s1_chipselect),                    //                                           .chipselect
		.ledOpcao3_s1_address                             (mm_interconnect_0_ledopcao3_s1_address),                       //                               ledOpcao3_s1.address
		.ledOpcao3_s1_write                               (mm_interconnect_0_ledopcao3_s1_write),                         //                                           .write
		.ledOpcao3_s1_readdata                            (mm_interconnect_0_ledopcao3_s1_readdata),                      //                                           .readdata
		.ledOpcao3_s1_writedata                           (mm_interconnect_0_ledopcao3_s1_writedata),                     //                                           .writedata
		.ledOpcao3_s1_chipselect                          (mm_interconnect_0_ledopcao3_s1_chipselect),                    //                                           .chipselect
		.ledOpcao4_s1_address                             (mm_interconnect_0_ledopcao4_s1_address),                       //                               ledOpcao4_s1.address
		.ledOpcao4_s1_write                               (mm_interconnect_0_ledopcao4_s1_write),                         //                                           .write
		.ledOpcao4_s1_readdata                            (mm_interconnect_0_ledopcao4_s1_readdata),                      //                                           .readdata
		.ledOpcao4_s1_writedata                           (mm_interconnect_0_ledopcao4_s1_writedata),                     //                                           .writedata
		.ledOpcao4_s1_chipselect                          (mm_interconnect_0_ledopcao4_s1_chipselect),                    //                                           .chipselect
		.ledOpcao5_s1_address                             (mm_interconnect_0_ledopcao5_s1_address),                       //                               ledOpcao5_s1.address
		.ledOpcao5_s1_write                               (mm_interconnect_0_ledopcao5_s1_write),                         //                                           .write
		.ledOpcao5_s1_readdata                            (mm_interconnect_0_ledopcao5_s1_readdata),                      //                                           .readdata
		.ledOpcao5_s1_writedata                           (mm_interconnect_0_ledopcao5_s1_writedata),                     //                                           .writedata
		.ledOpcao5_s1_chipselect                          (mm_interconnect_0_ledopcao5_s1_chipselect),                    //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken)                   //                                           .clken
	);

	projeto1_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
