// ProjetoSemInstruction.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ProjetoSemInstruction (
		input  wire       botaodescer_external_connection_export, // botaodescer_external_connection.export
		input  wire       botaoentrar_external_connection_export, // botaoentrar_external_connection.export
		input  wire       botaosubir_external_connection_export,  //  botaosubir_external_connection.export
		input  wire       botaovoltar_external_connection_export, // botaovoltar_external_connection.export
		input  wire       clk_clk,                                //                             clk.clk
		output wire       lcd_16207_0_external_RS,                //            lcd_16207_0_external.RS
		output wire       lcd_16207_0_external_RW,                //                                .RW
		inout  wire [7:0] lcd_16207_0_external_data,              //                                .data
		output wire       lcd_16207_0_external_E,                 //                                .E
		output wire       ledazul_external_connection_export,     //     ledazul_external_connection.export
		output wire       ledverde_external_connection_export,    //    ledverde_external_connection.export
		output wire       ledvermelho_external_connection_export, // ledvermelho_external_connection.export
		input  wire       reset_reset_n                           //                           reset.reset_n
	);

	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [17:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [17:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_readdata;         // lcd_16207_0:readdata -> mm_interconnect_0:lcd_16207_0_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_16207_0_control_slave_address;          // mm_interconnect_0:lcd_16207_0_control_slave_address -> lcd_16207_0:address
	wire         mm_interconnect_0_lcd_16207_0_control_slave_read;             // mm_interconnect_0:lcd_16207_0_control_slave_read -> lcd_16207_0:read
	wire         mm_interconnect_0_lcd_16207_0_control_slave_begintransfer;    // mm_interconnect_0:lcd_16207_0_control_slave_begintransfer -> lcd_16207_0:begintransfer
	wire         mm_interconnect_0_lcd_16207_0_control_slave_write;            // mm_interconnect_0:lcd_16207_0_control_slave_write -> lcd_16207_0:write
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_writedata;        // mm_interconnect_0:lcd_16207_0_control_slave_writedata -> lcd_16207_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_ledazul_s1_chipselect;                      // mm_interconnect_0:ledAzul_s1_chipselect -> ledAzul:chipselect
	wire  [31:0] mm_interconnect_0_ledazul_s1_readdata;                        // ledAzul:readdata -> mm_interconnect_0:ledAzul_s1_readdata
	wire   [1:0] mm_interconnect_0_ledazul_s1_address;                         // mm_interconnect_0:ledAzul_s1_address -> ledAzul:address
	wire         mm_interconnect_0_ledazul_s1_write;                           // mm_interconnect_0:ledAzul_s1_write -> ledAzul:write_n
	wire  [31:0] mm_interconnect_0_ledazul_s1_writedata;                       // mm_interconnect_0:ledAzul_s1_writedata -> ledAzul:writedata
	wire         mm_interconnect_0_ledverde_s1_chipselect;                     // mm_interconnect_0:ledVerde_s1_chipselect -> ledVerde:chipselect
	wire  [31:0] mm_interconnect_0_ledverde_s1_readdata;                       // ledVerde:readdata -> mm_interconnect_0:ledVerde_s1_readdata
	wire   [1:0] mm_interconnect_0_ledverde_s1_address;                        // mm_interconnect_0:ledVerde_s1_address -> ledVerde:address
	wire         mm_interconnect_0_ledverde_s1_write;                          // mm_interconnect_0:ledVerde_s1_write -> ledVerde:write_n
	wire  [31:0] mm_interconnect_0_ledverde_s1_writedata;                      // mm_interconnect_0:ledVerde_s1_writedata -> ledVerde:writedata
	wire         mm_interconnect_0_ledvermelho_s1_chipselect;                  // mm_interconnect_0:ledVermelho_s1_chipselect -> ledVermelho:chipselect
	wire  [31:0] mm_interconnect_0_ledvermelho_s1_readdata;                    // ledVermelho:readdata -> mm_interconnect_0:ledVermelho_s1_readdata
	wire   [1:0] mm_interconnect_0_ledvermelho_s1_address;                     // mm_interconnect_0:ledVermelho_s1_address -> ledVermelho:address
	wire         mm_interconnect_0_ledvermelho_s1_write;                       // mm_interconnect_0:ledVermelho_s1_write -> ledVermelho:write_n
	wire  [31:0] mm_interconnect_0_ledvermelho_s1_writedata;                   // mm_interconnect_0:ledVermelho_s1_writedata -> ledVermelho:writedata
	wire  [31:0] mm_interconnect_0_botaovoltar_s1_readdata;                    // botaoVoltar:readdata -> mm_interconnect_0:botaoVoltar_s1_readdata
	wire   [1:0] mm_interconnect_0_botaovoltar_s1_address;                     // mm_interconnect_0:botaoVoltar_s1_address -> botaoVoltar:address
	wire  [31:0] mm_interconnect_0_botaoentrar_s1_readdata;                    // botaoEntrar:readdata -> mm_interconnect_0:botaoEntrar_s1_readdata
	wire   [1:0] mm_interconnect_0_botaoentrar_s1_address;                     // mm_interconnect_0:botaoEntrar_s1_address -> botaoEntrar:address
	wire  [31:0] mm_interconnect_0_botaodescer_s1_readdata;                    // botaoDescer:readdata -> mm_interconnect_0:botaoDescer_s1_readdata
	wire   [1:0] mm_interconnect_0_botaodescer_s1_address;                     // mm_interconnect_0:botaoDescer_s1_address -> botaoDescer:address
	wire  [31:0] mm_interconnect_0_botaosubir_s1_readdata;                     // botaoSubir:readdata -> mm_interconnect_0:botaoSubir_s1_readdata
	wire   [1:0] mm_interconnect_0_botaosubir_s1_address;                      // mm_interconnect_0:botaoSubir_s1_address -> botaoSubir:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [botaoDescer:reset_n, botaoEntrar:reset_n, botaoSubir:reset_n, botaoVoltar:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, lcd_16207_0:reset_n, ledAzul:reset_n, ledVerde:reset_n, ledVermelho:reset_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	ProjetoSemInstruction_botaoDescer botaodescer (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_botaodescer_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botaodescer_s1_readdata), //                    .readdata
		.in_port  (botaodescer_external_connection_export)     // external_connection.export
	);

	ProjetoSemInstruction_botaoDescer botaoentrar (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_botaoentrar_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botaoentrar_s1_readdata), //                    .readdata
		.in_port  (botaoentrar_external_connection_export)     // external_connection.export
	);

	ProjetoSemInstruction_botaoDescer botaosubir (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_botaosubir_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botaosubir_s1_readdata), //                    .readdata
		.in_port  (botaosubir_external_connection_export)     // external_connection.export
	);

	ProjetoSemInstruction_botaoDescer botaovoltar (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_botaovoltar_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botaovoltar_s1_readdata), //                    .readdata
		.in_port  (botaovoltar_external_connection_export)     // external_connection.export
	);

	ProjetoSemInstruction_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	ProjetoSemInstruction_lcd_16207_0 lcd_16207_0 (
		.reset_n       (~rst_controller_reset_out_reset),                           //         reset.reset_n
		.clk           (clk_clk),                                                   //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_16207_0_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_16207_0_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_16207_0_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_16207_0_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_16207_0_control_slave_address),       //              .address
		.LCD_RS        (lcd_16207_0_external_RS),                                   //      external.export
		.LCD_RW        (lcd_16207_0_external_RW),                                   //              .export
		.LCD_data      (lcd_16207_0_external_data),                                 //              .export
		.LCD_E         (lcd_16207_0_external_E)                                     //              .export
	);

	ProjetoSemInstruction_ledAzul ledazul (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_ledazul_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledazul_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledazul_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledazul_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledazul_s1_readdata),   //                    .readdata
		.out_port   (ledazul_external_connection_export)       // external_connection.export
	);

	ProjetoSemInstruction_ledAzul ledverde (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_ledverde_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledverde_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledverde_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledverde_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledverde_s1_readdata),   //                    .readdata
		.out_port   (ledverde_external_connection_export)       // external_connection.export
	);

	ProjetoSemInstruction_ledAzul ledvermelho (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_ledvermelho_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledvermelho_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledvermelho_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledvermelho_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledvermelho_s1_readdata),   //                    .readdata
		.out_port   (ledvermelho_external_connection_export)       // external_connection.export
	);

	ProjetoSemInstruction_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	ProjetoSemInstruction_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	ProjetoSemInstruction_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.botaoDescer_s1_address                           (mm_interconnect_0_botaodescer_s1_address),                     //                             botaoDescer_s1.address
		.botaoDescer_s1_readdata                          (mm_interconnect_0_botaodescer_s1_readdata),                    //                                           .readdata
		.botaoEntrar_s1_address                           (mm_interconnect_0_botaoentrar_s1_address),                     //                             botaoEntrar_s1.address
		.botaoEntrar_s1_readdata                          (mm_interconnect_0_botaoentrar_s1_readdata),                    //                                           .readdata
		.botaoSubir_s1_address                            (mm_interconnect_0_botaosubir_s1_address),                      //                              botaoSubir_s1.address
		.botaoSubir_s1_readdata                           (mm_interconnect_0_botaosubir_s1_readdata),                     //                                           .readdata
		.botaoVoltar_s1_address                           (mm_interconnect_0_botaovoltar_s1_address),                     //                             botaoVoltar_s1.address
		.botaoVoltar_s1_readdata                          (mm_interconnect_0_botaovoltar_s1_readdata),                    //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.lcd_16207_0_control_slave_address                (mm_interconnect_0_lcd_16207_0_control_slave_address),          //                  lcd_16207_0_control_slave.address
		.lcd_16207_0_control_slave_write                  (mm_interconnect_0_lcd_16207_0_control_slave_write),            //                                           .write
		.lcd_16207_0_control_slave_read                   (mm_interconnect_0_lcd_16207_0_control_slave_read),             //                                           .read
		.lcd_16207_0_control_slave_readdata               (mm_interconnect_0_lcd_16207_0_control_slave_readdata),         //                                           .readdata
		.lcd_16207_0_control_slave_writedata              (mm_interconnect_0_lcd_16207_0_control_slave_writedata),        //                                           .writedata
		.lcd_16207_0_control_slave_begintransfer          (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer),    //                                           .begintransfer
		.ledAzul_s1_address                               (mm_interconnect_0_ledazul_s1_address),                         //                                 ledAzul_s1.address
		.ledAzul_s1_write                                 (mm_interconnect_0_ledazul_s1_write),                           //                                           .write
		.ledAzul_s1_readdata                              (mm_interconnect_0_ledazul_s1_readdata),                        //                                           .readdata
		.ledAzul_s1_writedata                             (mm_interconnect_0_ledazul_s1_writedata),                       //                                           .writedata
		.ledAzul_s1_chipselect                            (mm_interconnect_0_ledazul_s1_chipselect),                      //                                           .chipselect
		.ledVerde_s1_address                              (mm_interconnect_0_ledverde_s1_address),                        //                                ledVerde_s1.address
		.ledVerde_s1_write                                (mm_interconnect_0_ledverde_s1_write),                          //                                           .write
		.ledVerde_s1_readdata                             (mm_interconnect_0_ledverde_s1_readdata),                       //                                           .readdata
		.ledVerde_s1_writedata                            (mm_interconnect_0_ledverde_s1_writedata),                      //                                           .writedata
		.ledVerde_s1_chipselect                           (mm_interconnect_0_ledverde_s1_chipselect),                     //                                           .chipselect
		.ledVermelho_s1_address                           (mm_interconnect_0_ledvermelho_s1_address),                     //                             ledVermelho_s1.address
		.ledVermelho_s1_write                             (mm_interconnect_0_ledvermelho_s1_write),                       //                                           .write
		.ledVermelho_s1_readdata                          (mm_interconnect_0_ledvermelho_s1_readdata),                    //                                           .readdata
		.ledVermelho_s1_writedata                         (mm_interconnect_0_ledvermelho_s1_writedata),                   //                                           .writedata
		.ledVermelho_s1_chipselect                        (mm_interconnect_0_ledvermelho_s1_chipselect),                  //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken)                   //                                           .clken
	);

	ProjetoSemInstruction_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
